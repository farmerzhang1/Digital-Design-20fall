module three_tb();
    reg [7:0] a, b;
    wire [7:0] c, d, e, f, g, h, i, j, k;